module state_switch(
	input CLK, RESET, X,
	output [3:0] state_out);

	typedef enum logic[3:0] {
		A1 = 4'b0000,
		A2 = 4'b0100,
		A3 = 4'b0001,
		A4 = 4'b0110,
		A5 = 4'b1100,
		A6 = 4'b0011,
		A7 = 4'b1001,
		A8 = 4'b1000,
		A9 = 4'b0010,
		A10 = 4'b0101}
	statetype;

	statetype state, next_state;
	
	always_ff @(posedge CLK, posedge RESET)
		if (RESET) state <= A1;
		else state <= next_state;
	
	always_comb
		case (state)
			A1: next_state <= X ? A2 : A3;
			A2: next_state <= X ? A4 : A5;
			A3: next_state <= X ? A6 : A7;
			A4: next_state <= X ? A8 : A9;
			A5: next_state <= A8;
			A6: next_state <= A9;
			A7: next_state <= X ? A9 : A8;
			A8: next_state <= A1;
			A9: next_state <= X ? A1 : A10;
			A10: next_state <= X ? A2 : A3;
			default: next_state <= A1;
		endcase
	
	assign state_out = state;
	
endmodule


module user_sequence(
	input CLK, RESET, X,
	output [3:0] sequence_out, slots);

	logic [3:0] user_sequence, slots_;
	
	always_ff @(posedge CLK, posedge RESET)
		if (RESET) slots_ = 4'b0000;
		else
			if (slots_[3]) slots_[3:1] = 3'b000;
			else
				begin
					slots_ = slots_ << 1;
					slots_[0] = 1;
				end

	always_ff @(posedge CLK)
		begin
			user_sequence = user_sequence << 1;
			user_sequence[0] = X;
		end
	
	assign slots = slots_;
	assign sequence_out = user_sequence;

endmodule


module digits_tube(
	input CLK_50M,
	input [3:0] state, user_sequence, slots,
	output [7:0] dataout,
	output [7:0] bit_out);
	
	typedef enum logic[7:0]{
		D0 = 8'b1100_0000,
		D1 = 8'b1111_1001,
		DM = 8'b1011_1111
		}digit;
	
	typedef enum logic[7:0]{
		B1 = 8'b1111_1110,
		B2 = 8'b1111_1101,
		B3 = 8'b1111_1011,
		B4 = 8'b1111_0111,
		B5 = 8'b1110_1111,
		B6 = 8'b1101_1111,
		B7 = 8'b1011_1111,
		B8 = 8'b0111_1111
	}slot;

	digit dataout_;
	slot bit_out_;
	bit [15:0] count;
	
	always @(posedge CLK_50M)
		if (count == 16'b1111111111111111) count = 0;
		else count = count + 1;
	
	always_ff @(posedge count[15])
		if (bit_out_ == B8) bit_out_ = B1;
		else bit_out_ = bit_out_.next();
	
	always_comb
		case(bit_out_)
			B1: dataout_ = slots[0] ? (user_sequence[0] ? D1:D0) : DM;
			B2: dataout_ = slots[1] ? (user_sequence[1] ? D1:D0) : DM;
			B3: dataout_ = slots[2] ? (user_sequence[2] ? D1:D0) : DM;
			B4: dataout_ = slots[3] ? (user_sequence[3] ? D1:D0) : DM;
			B5: dataout_ = state[0] ? D1:D0;
			B6: dataout_ = state[1] ? D1:D0;
			B7: dataout_ = state[2] ? D1:D0;
			B8: dataout_ = state[3] ? D1:D0;
			default: dataout_ = D0;
		endcase
	
	assign dataout = dataout_;
	assign bit_out = bit_out_;

endmodule

module always_one(
	output one);
	
	assign one = 1;

endmodule


/*module state_machine_lab2(
	input RESET, X0, X1,
	input CLK_50M,
	output [11: 0] Y,
	output [7:0] dataout,
	output [7:0] bit_out);

	
	bit [3:0] A10 = 4'b0101;
	logic CLK_;
	logic [3:0] state, user_sequence, slots;
	
	assign CLK_ = X0 ^ X1;
	
	state_switch get_state(CLK_, RESET, X1, state);
	user_sequence get_sequence(CLK_, RESET, X1, user_sequence, slots);
	digits_tube display(CLK_50M, state, user_sequence, slots, dataout, bit_out);
	assign Y = {12{state == A10 & CLK_}};

endmodule*/
